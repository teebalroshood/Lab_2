
`default_nettype none

module circuit_A_v2(
	input 	i_v3,
	input 	i_v2,
	input 	i_v1,
	input 	i_v0,
	output 	o_a0,
	output 	o_a1,
	output 	o_a2,
	output 	o_a3
);

	// Combinational Logic only
	// TODO

endmodule
